`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:05:51 10/02/2015 
// Design Name: 
// Module Name:    traffic_light_hw 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module traffic_light_hw(
    input clk,
    input reset,
    output reg green_light , red_light, yellow_light,
	output reg [3:0] cnt 
    );



endmodule
